library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity aes is
generic
	(
		DATA_WIDTH_AES : natural := 128
	);
  port(
    msg : in std_logic_vector(0 to 127);
	 mensagem_criptografada : out std_logic_vector(0 to 63) ;
	 clk		  : in std_logic;
	 reset : in std_logic;
	 En_regAdder: in std_logic
  );
end aes;

architecture inst_aes of aes is
  type matriz is array (integer range 0 to 15) of std_logic_vector (0 to 7);
  type subByte is array (integer range 0 to 255) of std_logic_vector(0 to 7);
  signal State, Cipherkey : matriz;
  signal Key : std_logic_vector(0 to 127);
  signal TabSubBytes : subByte;
  signal temp : std_logic_vector(0 to 7);
  signal outMux1, outMux2, outAdder, outRegAdder, outRegA, outRegB, outInv : std_logic_vector  ((DATA_WIDTH_AES-1) downto 0);
  

component registerNbits is

	generic
	(
		DATA_WIDTH : natural := 128
	);

	port 
	(
		clk		: in std_logic;
		enable	: in std_logic;
		d	      : in std_logic_vector((DATA_WIDTH-1) downto 0);
		q			: out std_logic_vector((DATA_WIDTH-1) downto 0)
		
	);

end component;  
  
component PC_AES is
    PORT (
		  -- Portas principais
        reset : in std_logic;
        clock : in std_logic;
        en_inputs : out std_logic;
        cTRL_mux1 : out std_logic;
        cTRL_mux2 : out std_logic;
        en_regULA : out std_logic;
		  -- Portas para depuração
		  state_view : out std_logic_vector(2 downto 0)
    );
END component;  
  
begin 

PC: 	PC_AES
			 --generic map (DATA_WIDTH_AES => GLOBAL_DATA_WIDTH)
			 port map (
						-- Portas de depuração
							clock => clk,
							reset => reset
						--	a_PO => a_top,
					--		b_PO => b_top,
					--		Ctrl_mux1 => ctrl_mux1_conect,
					--		Ctrl_mux2 => Ctrl_mux2_conect,
						--	en_inputs => en_inputs_conect,
							--en_regAdder => en_regAdder_conect,
							--c_PO => c_top,
							
						-- Portas de depuração
					--		outMux1_view => outMux1_view,
						--	outMux2_view => outMux2_view, 
							--outAdder_view => outAdder_view, 
			--				outRegAdder_view => outRegAdder_view, 
				--			outRegA_view => outRegA_view, 
					--		outRegB_view => outRegB_view, 
						--	outInv_view => outInv_view
						);	
						
RegAdder: 	registerNbits
			 generic map (DATA_WIDTH => DATA_WIDTH_AES)
			 port map (clk => clk, enable => En_regAdder, d => outAdder, q => outRegAdder);	
  --          0000    0001    0002    0003    0004    0005    0006    0007    0008    0009    0000    0001    0002    0003    0004    0005                                                                                            
  Key <= "00110000001100010011001000110011001101000011010100110110001101110011100000111001001100000011000100110010001100110011010000110101";
  process(clk)
  --Declaração de variáveis
  variable posicao : integer;
  --variable temp : std_logic_vector(0 to 7);
  --Fim de declaração de variáveis
  begin 

    --Assinala a mensagem a ser criptografada na matriz state
	 for i in 0 to 15 loop 
      State(i) <= msg((120 - (i * 8)) to (127 - (i * 8)));
    end loop;
	 
    --Assinala a chave a ser utilizada(0123456789012345) na matriz key
	 for i in 0 to 15 loop 
      CipherKey(i) <= Key((120 - (i * 8)) to (127 - (i * 8)));
    end loop;
      
    --Faz o AddRoundKey
    for i in 0 to 15 loop 
	   for j in 0 to 7 loop 
        State(i)(j) <= State(i)(j) xor CipherKey(i)(j);
		end loop;  
    end loop;
	 
	
	 
	 --Etapa de SubBytes
	 for i in 0 to 15 loop 
	   posicao := to_integer(unsigned(State(i)(0 to 7)));
      State(i) <= TabSubBytes(posicao);
    end loop;
	 
	 --Etapa de ShiftRows
	 for i in 4 to 7 loop --Rotaciona um byte a esquerda
	 
	 end loop;
	 for i in 8 to 11 loop --Rotaciona duas vezes um byte a esquerda
	 
	 end loop;
	 for i in 12 to 15 loop --Rotaciona três vezes um byte a esquerda
	 
	 end loop;
	 
  end process;
  
end inst_aes;


