library ieee;
use ieee.std_logic_1164.all;

entity AddRoundKey is
 
end AddRoundKey;

architecture inst_AddRoundKey of AddRoundKey is
  type matriz is array (integer range 0 to 7) of std_logic_vector (15 downto 0);
  signal State, Cipherkey : matriz;

begin 
 
  
  
  
  
  
end inst_AddRoundKey;